`define HWDATA_WIDTH32
`define ADDR_WIDTH32
